`default_nettype none

module warp_hart (
    
);
    wire [63:0] buffer;
endmodule
