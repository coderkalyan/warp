`default_nettype none

// TODO: parametrize cache size
module warp_icache (
    input  wire [63:]
);
endmodule
